`timescale 1 ns/ 10 ps
module VT_RNG(data, data2, reset, clk, x);//V-trapezoid method Random Number Generator
input [38:0] data;
input [15:0] data2;
input  clk, reset;
output [17:0] x;

reg [38:0] lfsr;
reg [15:0] lfsr2;
reg [17:0] x;
reg [12:0] i_t0;
reg s,s_t1;
reg [3:0] mi,mi_t1,mi_t2;
reg [17:0] xl,xl_t1,xl_t2,xl_t3;
reg [12:0] ri,ri_t1;
reg [12:0] u1_t0,u2_t0,u3_t0,u1_t1,u2_t1,u3_t1;
reg q1,q1_t1;
reg [12:0] q2,q3,q3_t2;
reg [17:0] q4,q4_t3;


wire linear_feedback;
wire linear_feedback2;

//==================================================================================

assign linear_feedback = (lfsr[0]^lfsr[4]);
assign linear_feedback2 = (lfsr2[0] ^ lfsr2[2] ^ lfsr2[3] ^ lfsr2[5]);

// Time 0 --------------------------------------------------------------------------

always @(posedge clk  or negedge reset)
if (!reset) begin
  lfsr  <= data ;
  lfsr2 <= data2 ;
end else begin
lfsr	<= {linear_feedback, lfsr[38:1]};
lfsr2	<= {linear_feedback2, lfsr2[15:1]};
u1_t0	<= {lfsr[13:12],lfsr[1:0],lfsr[7:6],lfsr[21:20],lfsr[31:30],lfsr[27:26],lfsr[34]};
u2_t0	<= {lfsr[9:8],lfsr[23:22],lfsr[5:4],lfsr[17:16],lfsr[25:24],lfsr[37:36],lfsr[27]};
u3_t0	<= {lfsr[19:18],lfsr[3:2],lfsr[11:10],lfsr[15:14],lfsr[33:32],lfsr[29:28],lfsr[35]};
i_t0	<= {lfsr2[9:8],lfsr2[11:10],lfsr2[5:4],lfsr2[15:14],lfsr2[3:2],lfsr2[1:0],lfsr2[7]};
end

// Time 1 --------------------------------------------------------------------------

always @(*) begin
	if(i_t0 >= 13'b0000000000000 && i_t0 <= 13'b0000000001100) begin s = 1'b1; mi = 4'b1101; xl = 18'b00000_0001000000000; ri = 13'b1110011001111; end
	else if(i_t0 >= 13'b0000000001101 && i_t0 <= 13'b0000000100010) begin s = 1'b1; mi = 4'b1100; xl = 18'b00000_0001100000000; ri = 13'b1110000000100; end
	else if(i_t0 >= 13'b0000000100011 && i_t0 <= 13'b0000000110011) begin s = 1'b1; mi = 4'b1100; xl = 18'b00000_0010100000000; ri = 13'b1110101100101; end
	else if(i_t0 >= 13'b0000000110100 && i_t0 <= 13'b0000001010001) begin s = 1'b1; mi = 4'b1011; xl = 18'b00000_0011100000000; ri = 13'b1110010010000; end
	else if(i_t0 >= 13'b0000001010010 && i_t0 <= 13'b0000001101001) begin s = 1'b1; mi = 4'b1011; xl = 18'b00000_0101100000000; ri = 13'b1110110110011; end
	else if(i_t0 >= 13'b0000001101010 && i_t0 <= 13'b0000010010010) begin s = 1'b1; mi = 4'b1010; xl = 18'b00000_0111100000000; ri = 13'b1110011111101; end
	else if(i_t0 >= 13'b0000010010011 && i_t0 <= 13'b0000010110101) begin s = 1'b1; mi = 4'b1010; xl = 18'b00000_1011100000000; ri = 13'b1111000011001; end
	else if(i_t0 >= 13'b0000010110110 && i_t0 <= 13'b0000011110100) begin s = 1'b1; mi = 4'b1001; xl = 18'b00000_1111100000000; ri = 13'b1110111111000; end
	else if(i_t0 >= 13'b0000011110101 && i_t0 <= 13'b0000100101101) begin s = 1'b1; mi = 4'b1001; xl = 18'b00001_0111100000000; ri = 13'b1111110000001; end
	else if(i_t0 >= 13'b0000100101110 && i_t0 <= 13'b0000101100111) begin s = 1'b0; mi = 4'b1001; xl = 18'b00001_1111100000000; ri = 13'b1111101010010; end
	else if(i_t0 >= 13'b0000101101000 && i_t0 <= 13'b0000110100110) begin s = 1'b0; mi = 4'b1001; xl = 18'b00010_0111100000000; ri = 13'b1111001011001; end
	else if(i_t0 >= 13'b0000110100111 && i_t0 <= 13'b0000111101101) begin s = 1'b0; mi = 4'b1001; xl = 18'b00010_1111100000000; ri = 13'b1110110010101; end
	else if(i_t0 >= 13'b0000111101110 && i_t0 <= 13'b0001001000001) begin s = 1'b0; mi = 4'b1001; xl = 18'b00011_0111100000000; ri = 13'b1110100001100; end
	else if(i_t0 >= 13'b0001001000010 && i_t0 <= 13'b0001010100111) begin s = 1'b0; mi = 4'b1001; xl = 18'b00011_1111100000000; ri = 13'b1110010111110; end
	else if(i_t0 >= 13'b0001010101000 && i_t0 <= 13'b0001100100101) begin s = 1'b0; mi = 4'b1001; xl = 18'b00100_0111100000000; ri = 13'b1110010100011; end
	else if(i_t0 >= 13'b0001100100110 && i_t0 <= 13'b0001110111111) begin s = 1'b0; mi = 4'b1001; xl = 18'b00100_1111100000000; ri = 13'b1110010110001; end
	else if(i_t0 >= 13'b0001111000000 && i_t0 <= 13'b0010001111101) begin s = 1'b0; mi = 4'b1001; xl = 18'b00101_0111100000000; ri = 13'b1110011011100; end
	else if(i_t0 >= 13'b0010001111110 && i_t0 <= 13'b0011001110010) begin s = 1'b0; mi = 4'b0000; xl = 18'b00101_1111100000000; ri = 13'b1101010010011; end
	else if(i_t0 >= 13'b0011001110011 && i_t0 <= 13'b0100100010010) begin s = 1'b0; mi = 4'b0000; xl = 18'b00110_1111100000000; ri = 13'b1101111101101; end
	else if(i_t0 >= 13'b0100100010011 && i_t0 <= 13'b0101010011111) begin s = 1'b0; mi = 4'b1001; xl = 18'b00111_1111100000000; ri = 13'b1111010001001; end
	else if(i_t0 >= 13'b0101010100000 && i_t0 <= 13'b0110001001100) begin s = 1'b0; mi = 4'b1001; xl = 18'b01000_0111100000000; ri = 13'b1111011110000; end
	else if(i_t0 >= 13'b0110001001101 && i_t0 <= 13'b0111000010000) begin s = 1'b0; mi = 4'b1001; xl = 18'b01000_1111100000000; ri = 13'b1111101011001; end
	else if(i_t0 >= 13'b0111000010001 && i_t0 <= 13'b0111111100001) begin s = 1'b0; mi = 4'b1001; xl = 18'b01001_0111100000000; ri = 13'b1111111000011; end
	else if(i_t0 >= 13'b0111111100010 && i_t0 <= 13'b1000110110011) begin s = 1'b1; mi = 4'b1001; xl = 18'b01001_1111100000000; ri = 13'b1111111010001; end
	else if(i_t0 >= 13'b1000110110100 && i_t0 <= 13'b1001101111010) begin s = 1'b1; mi = 4'b1001; xl = 18'b01010_0111100000000; ri = 13'b1111101100110; end
	else if(i_t0 >= 13'b1001101111011 && i_t0 <= 13'b1010100101010) begin s = 1'b1; mi = 4'b1001; xl = 18'b01010_1111100000000; ri = 13'b1111011111101; end
	else if(i_t0 >= 13'b1010100101011 && i_t0 <= 13'b1011010111100) begin s = 1'b1; mi = 4'b1001; xl = 18'b01011_0111100000000; ri = 13'b1111010010101; end
	else if(i_t0 >= 13'b1011010111101 && i_t0 <= 13'b1100101100110) begin s = 1'b1; mi = 4'b0000; xl = 18'b01011_1111100000000; ri = 13'b1110000000101; end
	else if(i_t0 >= 13'b1100101100111 && i_t0 <= 13'b1101101100101) begin s = 1'b1; mi = 4'b0000; xl = 18'b01100_1111100000000; ri = 13'b1101010100110; end
	else if(i_t0 >= 13'b1101101100110 && i_t0 <= 13'b1110000101000) begin s = 1'b1; mi = 4'b1001; xl = 18'b01101_1111100000000; ri = 13'b1110011100011; end
	else if(i_t0 >= 13'b1110000101001 && i_t0 <= 13'b1110011000111) begin s = 1'b1; mi = 4'b1001; xl = 18'b01110_0111100000000; ri = 13'b1110010110101; end
	else if(i_t0 >= 13'b1110011001000 && i_t0 <= 13'b1110101001000) begin s = 1'b1; mi = 4'b1001; xl = 18'b01110_1111100000000; ri = 13'b1110010100011; end
	else if(i_t0 >= 13'b1110101001001 && i_t0 <= 13'b1110110110001) begin s = 1'b1; mi = 4'b1001; xl = 18'b01111_0111100000000; ri = 13'b1110010111000; end
	else if(i_t0 >= 13'b1110110110010 && i_t0 <= 13'b1111000000111) begin s = 1'b1; mi = 4'b1001; xl = 18'b01111_1111100000000; ri = 13'b1110011111111; end
	else if(i_t0 >= 13'b1111000001000 && i_t0 <= 13'b1111001001111) begin s = 1'b1; mi = 4'b1001; xl = 18'b10000_0111100000000; ri = 13'b1110110000001; end
	else if(i_t0 >= 13'b1111001010000 && i_t0 <= 13'b1111010001110) begin s = 1'b1; mi = 4'b1001; xl = 18'b10000_1111100000000; ri = 13'b1111000111110; end
	else if(i_t0 >= 13'b1111010001111 && i_t0 <= 13'b1111011001000) begin s = 1'b1; mi = 4'b1001; xl = 18'b10001_0111100000000; ri = 13'b1111100110000; end
	else if(i_t0 >= 13'b1111011001001 && i_t0 <= 13'b1111100000010) begin s = 1'b0; mi = 4'b1001; xl = 18'b10001_1111100000000; ri = 13'b1111110101010; end
	else if(i_t0 >= 13'b1111100000011 && i_t0 <= 13'b1111100111111) begin s = 1'b0; mi = 4'b1001; xl = 18'b10010_0111100000000; ri = 13'b1111000110011; end
	else if(i_t0 >= 13'b1111101000000 && i_t0 <= 13'b1111101100001) begin s = 1'b0; mi = 4'b1010; xl = 18'b10010_1111100000000; ri = 13'b1111001001010; end
	else if(i_t0 >= 13'b1111101100010 && i_t0 <= 13'b1111110001001) begin s = 1'b0; mi = 4'b1010; xl = 18'b10011_0011100000000; ri = 13'b1110101010111; end
	else if(i_t0 >= 13'b1111110001010 && i_t0 <= 13'b1111110011111) begin s = 1'b0; mi = 4'b1011; xl = 18'b10011_0111100000000; ri = 13'b1111000001010; end
	else if(i_t0 >= 13'b1111110100000 && i_t0 <= 13'b1111110111010) begin s = 1'b0; mi = 4'b1011; xl = 18'b10011_1001100000000; ri = 13'b1110100111100; end
	else if(i_t0 >= 13'b1111110111011 && i_t0 <= 13'b1111111011011) begin s = 1'b0; mi = 4'b1011; xl = 18'b10011_1011100000000; ri = 13'b1101101111101; end
	else if(i_t0 >= 13'b1111111011100 && i_t0 <= 13'b1111111110001) begin s = 1'b0; mi = 4'b1100; xl = 18'b10011_1101100000000; ri = 13'b1110000000100; end
	else if(i_t0 >= 13'b1111111110010 && i_t0 <= 13'b1111111111111) begin s = 1'b0; mi = 4'b1101; xl = 18'b10011_1110100000000; ri = 13'b1110011001111; end

	if(u2_t0 < u3_t0) begin q1 = 1; end
	else if(u2_t0 > u3_t0) begin q1 = 0;end
end

always @(posedge clk)
begin
	s_t1 <= s;
	mi_t1 <= mi;
	xl_t1 <= xl;
	ri_t1 <= ri;
	u1_t1 <= u1_t0;
	u2_t1 <= u2_t0;
	u3_t1 <= u3_t0;
	q1_t1 <= q1;
end

// Time 2 --------------------------------------------------------------------------

always @(*) begin
	q2 = (s_t1 ^ q1_t1) ? u3_t1 : u2_t1;
	q3 = (u1_t1 < ri_t1) ? u2_t1 : q2;
end

always @(posedge clk)
begin
	q3_t2 <= q3;
	mi_t2 <= mi_t1;
	xl_t2 <= xl_t1;
end


// Time 3 --------------------------------------------------------------------------

always @(*) begin
	q4 = (mi_t2[3]) ? q3_t2 >> mi_t2[2:0] : q3_t2 << mi_t2[2:0];
end

always @(posedge clk)
begin
	xl_t3 <= xl_t2;
	q4_t3 <= q4;
end

// Time 4 --------------------------------------------------------------------------

always @(posedge clk)
begin
	x <= q4_t3 + xl_t3;
end

//==================================================================================

endmodule
